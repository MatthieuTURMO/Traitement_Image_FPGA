----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:30:16 11/16/2015 
-- Design Name: 
-- Module Name:    Basc_D_1b - Basc_D_1b_arch 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Basc_D_1b is
    Port ( RESET : in STD_LOGIC;
           CLK : in  STD_LOGIC;
			   D : in  STD_LOGIC;
           Q : out  STD_LOGIC);
end Basc_D_1b;

architecture Basc_D_1b_arch of Basc_D_1b is

begin

process(CLK)
begin

if(RESET = '0') then
	if(CLK'event and CLK = '1') then
		Q<=D;
	end if;
else
		Q <= '0';
end if;
end process;



end Basc_D_1b_arch;

